`timescale 1ns / 1ps
//d1 approximation
module adder_tree_De2AXA( input wire [7:0]a,b,c,d,e,f,g,h, 
                    input wire clk, rst,
                   output wire [10:0]y );

reg [8:0] i11,i12,i13,i14;
reg [9:0] i21, i22;
reg [10:0] i31;
reg itest;
always@(posedge clk, posedge rst) begin
 if(rst) begin
 i11<=0; 
 i12<=0; 
 i13<=0; 
 i14<=0; 
 i21<=0;
 i31<=0;


 end
 else begin
 i11<= {a[7:3]+b[7:3]+(a[2]*b[2]) , ((a[2]*b[2])? 1'b0 : (a[2]+b[2])) + a[1]*b[1] ,a[1]+b[1], 1'b1};
 i12<= {c[7:3]+d[7:3]+(c[2]*d[2]) , ((c[2]*d[2])? 1'b0 : (c[2]+d[2])) + c[1]*d[1] ,c[1]+d[1], 1'b1};
 i13<= {e[7:3]+f[7:3]+(e[2]*f[2]) , ((e[2]*f[2])? 1'b0 : (e[2]+f[2])) + e[1]*f[1] ,e[1]+f[1], 1'b1};
 i14<= {g[7:3]+h[7:3]+(g[2]*h[2]) , ((g[2]*h[2])? 1'b0 : (g[2]+h[2])) + g[1]*h[1],g[1]+h[1], 1'b1};
 i21<= {i11[8:3]+i12[8:3]+(i11[2]*i12[2]), ((i11[2]*i12[2])? 1'b0 : (i11[2]+i12[2])) + i11[1]*i12[1] ,i11[1]+i12[1], 1'b1};
 i22<= {i13[8:3]+i14[8:3]+(i13[2]*i14[2]), ((i13[2]*i14[2])? 1'b0 : (i13[2]+i14[2])) + i13[1]*i14[1] ,i13[1]+i14[1], 1'b1};
 i31<= {i21[9:3]+i22[9:3]+(i21[2]*i22[2]), ((i21[2]*i22[2])? 1'b0 : (i21[2]+i22[2])) + i21[1]*i22[1] ,i21[1]+i22[1], 1'b1};

 end
 
end 


assign y = i31;


endmodule
